// BINARY TO BCD
module BIN2BCD	( 
// 
);


endmodule
