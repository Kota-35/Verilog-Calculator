// BCD TO BINARY
module BCD2BIN	( 
// 
);


endmodule
